// RTL (Verilog) generated @ Sat Mar 14 23:52:48 2020 by V3 
//               compiled @ Mar  7 2020 15:04:17
// Internal nets are renamed with prefix "v3_1584201168_".

// Module vendingMachine
module vendingMachine
(
   clk,
   reset,
   coinInNTD_50,
   coinInNTD_10,
   coinInNTD_5,
   coinInNTD_1,
   itemTypeIn,
   p,
   coinOutNTD_50,
   coinOutNTD_10,
   coinOutNTD_5,
   coinOutNTD_1,
   itemTypeOut,
   serviceTypeOut
);

   // Clock Signal for Synchronous DFF
   input clk;

   // I/O Declarations
   input reset;
   input [1:0] coinInNTD_50;
   input [1:0] coinInNTD_10;
   input [1:0] coinInNTD_5;
   input [1:0] coinInNTD_1;
   input [1:0] itemTypeIn;
   output p;
   output [2:0] coinOutNTD_50;
   output [2:0] coinOutNTD_10;
   output [2:0] coinOutNTD_5;
   output [2:0] coinOutNTD_1;
   output [1:0] itemTypeOut;
   output [1:0] serviceTypeOut;

   // Wire and Reg Declarations
   wire v3_1584201168_0;
   wire clk;
   wire reset;
   wire [1:0] coinInNTD_50;
   wire [1:0] coinInNTD_10;
   wire [1:0] coinInNTD_5;
   wire [1:0] coinInNTD_1;
   wire [1:0] itemTypeIn;
   reg [2:0] v3_1584201168_8;
   reg [2:0] v3_1584201168_9;
   reg [2:0] v3_1584201168_10;
   reg [2:0] v3_1584201168_11;
   reg [1:0] v3_1584201168_12;
   reg [1:0] v3_1584201168_13;
   reg v3_1584201168_14;
   reg [7:0] v3_1584201168_15;
   reg v3_1584201168_16;
   reg [1:0] v3_1584201168_17;
   reg [7:0] v3_1584201168_18;
   reg [2:0] v3_1584201168_19;
   reg [2:0] v3_1584201168_20;
   reg [2:0] v3_1584201168_21;
   reg [2:0] v3_1584201168_22;
   wire [2:0] v3_1584201168_23;
   wire [2:0] v3_1584201168_24;
   wire [2:0] v3_1584201168_25;
   wire [2:0] v3_1584201168_26;
   wire [2:0] v3_1584201168_27;
   wire [2:0] v3_1584201168_28;
   wire [2:0] v3_1584201168_29;
   wire [2:0] v3_1584201168_30;
   wire [2:0] v3_1584201168_31;
   wire [2:0] v3_1584201168_32;
   wire [2:0] v3_1584201168_33;
   wire [2:0] v3_1584201168_34;
   wire [2:0] v3_1584201168_35;
   wire v3_1584201168_36;
   wire v3_1584201168_37;
   wire [7:0] v3_1584201168_38;
   wire v3_1584201168_39;
   wire [1:0] v3_1584201168_40;
   wire v3_1584201168_41;
   wire [1:0] v3_1584201168_42;
   wire [2:0] v3_1584201168_43;
   wire [2:0] v3_1584201168_44;
   wire [2:0] v3_1584201168_45;
   wire [2:0] v3_1584201168_46;
   wire [2:0] v3_1584201168_47;
   wire v3_1584201168_48;
   wire v3_1584201168_49;
   wire [7:0] v3_1584201168_50;
   wire v3_1584201168_51;
   wire [1:0] v3_1584201168_52;
   wire v3_1584201168_53;
   wire [2:0] v3_1584201168_54;
   wire v3_1584201168_55;
   wire [2:0] v3_1584201168_56;
   wire [2:0] v3_1584201168_57;
   wire v3_1584201168_58;
   wire v3_1584201168_59;
   wire v3_1584201168_60;
   wire [2:0] v3_1584201168_61;
   wire v3_1584201168_62;
   wire [2:0] v3_1584201168_63;
   wire [2:0] v3_1584201168_64;
   wire [2:0] v3_1584201168_65;
   wire [2:0] v3_1584201168_66;
   wire [2:0] v3_1584201168_67;
   wire [2:0] v3_1584201168_68;
   wire [2:0] v3_1584201168_69;
   wire [2:0] v3_1584201168_70;
   wire [2:0] v3_1584201168_71;
   wire [2:0] v3_1584201168_72;
   wire [2:0] v3_1584201168_73;
   wire [2:0] v3_1584201168_74;
   wire [2:0] v3_1584201168_75;
   wire [2:0] v3_1584201168_76;
   wire [2:0] v3_1584201168_77;
   wire [2:0] v3_1584201168_78;
   wire [2:0] v3_1584201168_79;
   wire v3_1584201168_80;
   wire v3_1584201168_81;
   wire [7:0] v3_1584201168_82;
   wire [2:0] v3_1584201168_83;
   wire [2:0] v3_1584201168_84;
   wire [2:0] v3_1584201168_85;
   wire [2:0] v3_1584201168_86;
   wire [2:0] v3_1584201168_87;
   wire [2:0] v3_1584201168_88;
   wire [2:0] v3_1584201168_89;
   wire [2:0] v3_1584201168_90;
   wire [2:0] v3_1584201168_91;
   wire [2:0] v3_1584201168_92;
   wire [2:0] v3_1584201168_93;
   wire [2:0] v3_1584201168_94;
   wire [2:0] v3_1584201168_95;
   wire [2:0] v3_1584201168_96;
   wire [2:0] v3_1584201168_97;
   wire [2:0] v3_1584201168_98;
   wire [2:0] v3_1584201168_99;
   wire [2:0] v3_1584201168_100;
   wire [2:0] v3_1584201168_101;
   wire [2:0] v3_1584201168_102;
   wire [2:0] v3_1584201168_103;
   wire v3_1584201168_104;
   wire v3_1584201168_105;
   wire [7:0] v3_1584201168_106;
   wire [2:0] v3_1584201168_107;
   wire [2:0] v3_1584201168_108;
   wire [2:0] v3_1584201168_109;
   wire [2:0] v3_1584201168_110;
   wire [2:0] v3_1584201168_111;
   wire [2:0] v3_1584201168_112;
   wire [2:0] v3_1584201168_113;
   wire [2:0] v3_1584201168_114;
   wire [2:0] v3_1584201168_115;
   wire [2:0] v3_1584201168_116;
   wire [2:0] v3_1584201168_117;
   wire [2:0] v3_1584201168_118;
   wire [2:0] v3_1584201168_119;
   wire [2:0] v3_1584201168_120;
   wire [2:0] v3_1584201168_121;
   wire [2:0] v3_1584201168_122;
   wire [2:0] v3_1584201168_123;
   wire [2:0] v3_1584201168_124;
   wire [2:0] v3_1584201168_125;
   wire [2:0] v3_1584201168_126;
   wire [2:0] v3_1584201168_127;
   wire [2:0] v3_1584201168_128;
   wire [2:0] v3_1584201168_129;
   wire [2:0] v3_1584201168_130;
   wire [1:0] v3_1584201168_131;
   wire [1:0] v3_1584201168_132;
   wire [1:0] v3_1584201168_133;
   wire [1:0] v3_1584201168_134;
   wire [1:0] v3_1584201168_135;
   wire [1:0] v3_1584201168_136;
   wire [1:0] v3_1584201168_137;
   wire [1:0] v3_1584201168_138;
   wire [1:0] v3_1584201168_139;
   wire [1:0] v3_1584201168_140;
   wire [1:0] v3_1584201168_141;
   wire [1:0] v3_1584201168_142;
   wire [1:0] v3_1584201168_143;
   wire [1:0] v3_1584201168_144;
   wire v3_1584201168_145;
   wire v3_1584201168_146;
   wire [1:0] v3_1584201168_147;
   wire [1:0] v3_1584201168_148;
   wire [1:0] v3_1584201168_149;
   wire [1:0] v3_1584201168_150;
   wire [1:0] v3_1584201168_151;
   wire [1:0] v3_1584201168_152;
   wire [1:0] v3_1584201168_153;
   wire [1:0] v3_1584201168_154;
   wire [1:0] v3_1584201168_155;
   wire [1:0] v3_1584201168_156;
   wire [1:0] v3_1584201168_157;
   wire [1:0] v3_1584201168_158;
   wire [1:0] v3_1584201168_159;
   wire [1:0] v3_1584201168_160;
   wire [1:0] v3_1584201168_161;
   wire [1:0] v3_1584201168_162;
   wire [1:0] v3_1584201168_163;
   wire [1:0] v3_1584201168_164;
   wire [1:0] v3_1584201168_165;
   wire [1:0] v3_1584201168_166;
   wire [1:0] v3_1584201168_167;
   wire [1:0] v3_1584201168_168;
   wire [1:0] v3_1584201168_169;
   wire v3_1584201168_170;
   wire v3_1584201168_171;
   wire v3_1584201168_172;
   wire v3_1584201168_173;
   wire v3_1584201168_174;
   wire [7:0] v3_1584201168_175;
   wire [7:0] v3_1584201168_176;
   wire [7:0] v3_1584201168_177;
   wire [7:0] v3_1584201168_178;
   wire [7:0] v3_1584201168_179;
   wire [7:0] v3_1584201168_180;
   wire [7:0] v3_1584201168_181;
   wire [7:0] v3_1584201168_182;
   wire [7:0] v3_1584201168_183;
   wire [7:0] v3_1584201168_184;
   wire [5:0] v3_1584201168_185;
   wire [7:0] v3_1584201168_186;
   wire [7:0] v3_1584201168_187;
   wire [7:0] v3_1584201168_188;
   wire [7:0] v3_1584201168_189;
   wire [7:0] v3_1584201168_190;
   wire [7:0] v3_1584201168_191;
   wire [7:0] v3_1584201168_192;
   wire [7:0] v3_1584201168_193;
   wire [7:0] v3_1584201168_194;
   wire [7:0] v3_1584201168_195;
   wire [7:0] v3_1584201168_196;
   wire [7:0] v3_1584201168_197;
   wire [7:0] v3_1584201168_198;
   wire [7:0] v3_1584201168_199;
   wire [7:0] v3_1584201168_200;
   wire [7:0] v3_1584201168_201;
   wire [7:0] v3_1584201168_202;
   wire [7:0] v3_1584201168_203;
   wire [7:0] v3_1584201168_204;
   wire [7:0] v3_1584201168_205;
   wire v3_1584201168_206;
   wire v3_1584201168_207;
   wire v3_1584201168_208;
   wire v3_1584201168_209;
   wire v3_1584201168_210;
   wire v3_1584201168_211;
   wire v3_1584201168_212;
   wire v3_1584201168_213;
   wire v3_1584201168_214;
   wire v3_1584201168_215;
   wire v3_1584201168_216;
   wire v3_1584201168_217;
   wire v3_1584201168_218;
   wire v3_1584201168_219;
   wire [1:0] v3_1584201168_220;
   wire [1:0] v3_1584201168_221;
   wire [1:0] v3_1584201168_222;
   wire [1:0] v3_1584201168_223;
   wire [1:0] v3_1584201168_224;
   wire [1:0] v3_1584201168_225;
   wire [1:0] v3_1584201168_226;
   wire [1:0] v3_1584201168_227;
   wire [1:0] v3_1584201168_228;
   wire [1:0] v3_1584201168_229;
   wire [1:0] v3_1584201168_230;
   wire [1:0] v3_1584201168_231;
   wire [1:0] v3_1584201168_232;
   wire [1:0] v3_1584201168_233;
   wire [1:0] v3_1584201168_234;
   wire [1:0] v3_1584201168_235;
   wire [1:0] v3_1584201168_236;
   wire [1:0] v3_1584201168_237;
   wire [1:0] v3_1584201168_238;
   wire [1:0] v3_1584201168_239;
   wire [1:0] v3_1584201168_240;
   wire [1:0] v3_1584201168_241;
   wire [1:0] v3_1584201168_242;
   wire [1:0] v3_1584201168_243;
   wire [1:0] v3_1584201168_244;
   wire [1:0] v3_1584201168_245;
   wire [1:0] v3_1584201168_246;
   wire [1:0] v3_1584201168_247;
   wire [1:0] v3_1584201168_248;
   wire [7:0] v3_1584201168_249;
   wire [7:0] v3_1584201168_250;
   wire [7:0] v3_1584201168_251;
   wire [7:0] v3_1584201168_252;
   wire [7:0] v3_1584201168_253;
   wire [7:0] v3_1584201168_254;
   wire [7:0] v3_1584201168_255;
   wire [7:0] v3_1584201168_256;
   wire [7:0] v3_1584201168_257;
   wire [7:0] v3_1584201168_258;
   wire [7:0] v3_1584201168_259;
   wire [7:0] v3_1584201168_260;
   wire [7:0] v3_1584201168_261;
   wire [7:0] v3_1584201168_262;
   wire [7:0] v3_1584201168_263;
   wire [7:0] v3_1584201168_264;
   wire [7:0] v3_1584201168_265;
   wire [7:0] v3_1584201168_266;
   wire [7:0] v3_1584201168_267;
   wire [7:0] v3_1584201168_268;
   wire [7:0] v3_1584201168_269;
   wire [7:0] v3_1584201168_270;
   wire [7:0] v3_1584201168_271;
   wire [7:0] v3_1584201168_272;
   wire [7:0] v3_1584201168_273;
   wire [7:0] v3_1584201168_274;
   wire [7:0] v3_1584201168_275;
   wire [7:0] v3_1584201168_276;
   wire [7:0] v3_1584201168_277;
   wire [7:0] v3_1584201168_278;
   wire [7:0] v3_1584201168_279;
   wire [7:0] v3_1584201168_280;
   wire [7:0] v3_1584201168_281;
   wire [7:0] v3_1584201168_282;
   wire [7:0] v3_1584201168_283;
   wire v3_1584201168_284;
   wire [7:0] v3_1584201168_285;
   wire v3_1584201168_286;
   wire [7:0] v3_1584201168_287;
   wire v3_1584201168_288;
   wire [7:0] v3_1584201168_289;
   wire [7:0] v3_1584201168_290;
   wire [2:0] v3_1584201168_291;
   wire [2:0] v3_1584201168_292;
   wire [2:0] v3_1584201168_293;
   wire [2:0] v3_1584201168_294;
   wire [2:0] v3_1584201168_295;
   wire [2:0] v3_1584201168_296;
   wire [2:0] v3_1584201168_297;
   wire [2:0] v3_1584201168_298;
   wire [2:0] v3_1584201168_299;
   wire [2:0] v3_1584201168_300;
   wire [2:0] v3_1584201168_301;
   wire [2:0] v3_1584201168_302;
   wire [2:0] v3_1584201168_303;
   wire [2:0] v3_1584201168_304;
   wire [2:0] v3_1584201168_305;
   wire [2:0] v3_1584201168_306;
   wire [2:0] v3_1584201168_307;
   wire [2:0] v3_1584201168_308;
   wire [2:0] v3_1584201168_309;
   wire [2:0] v3_1584201168_310;
   wire [2:0] v3_1584201168_311;
   wire [2:0] v3_1584201168_312;
   wire [2:0] v3_1584201168_313;
   wire [2:0] v3_1584201168_314;
   wire v3_1584201168_315;
   wire [3:0] v3_1584201168_316;
   wire [3:0] v3_1584201168_317;
   wire [3:0] v3_1584201168_318;
   wire [3:0] v3_1584201168_319;
   wire [3:0] v3_1584201168_320;
   wire [3:0] v3_1584201168_321;
   wire [3:0] v3_1584201168_322;
   wire [2:0] v3_1584201168_323;
   wire [2:0] v3_1584201168_324;
   wire [2:0] v3_1584201168_325;
   wire [2:0] v3_1584201168_326;
   wire [2:0] v3_1584201168_327;
   wire [2:0] v3_1584201168_328;
   wire [2:0] v3_1584201168_329;
   wire [2:0] v3_1584201168_330;
   wire [2:0] v3_1584201168_331;
   wire [2:0] v3_1584201168_332;
   wire [2:0] v3_1584201168_333;
   wire [2:0] v3_1584201168_334;
   wire [2:0] v3_1584201168_335;
   wire [2:0] v3_1584201168_336;
   wire [2:0] v3_1584201168_337;
   wire [2:0] v3_1584201168_338;
   wire [2:0] v3_1584201168_339;
   wire [2:0] v3_1584201168_340;
   wire [2:0] v3_1584201168_341;
   wire [2:0] v3_1584201168_342;
   wire [2:0] v3_1584201168_343;
   wire [2:0] v3_1584201168_344;
   wire [2:0] v3_1584201168_345;
   wire [2:0] v3_1584201168_346;
   wire [2:0] v3_1584201168_347;
   wire [2:0] v3_1584201168_348;
   wire v3_1584201168_349;
   wire [3:0] v3_1584201168_350;
   wire [3:0] v3_1584201168_351;
   wire [3:0] v3_1584201168_352;
   wire [3:0] v3_1584201168_353;
   wire [3:0] v3_1584201168_354;
   wire [3:0] v3_1584201168_355;
   wire [2:0] v3_1584201168_356;
   wire [2:0] v3_1584201168_357;
   wire [2:0] v3_1584201168_358;
   wire [2:0] v3_1584201168_359;
   wire [2:0] v3_1584201168_360;
   wire [2:0] v3_1584201168_361;
   wire [2:0] v3_1584201168_362;
   wire [2:0] v3_1584201168_363;
   wire [2:0] v3_1584201168_364;
   wire [2:0] v3_1584201168_365;
   wire [2:0] v3_1584201168_366;
   wire [2:0] v3_1584201168_367;
   wire [2:0] v3_1584201168_368;
   wire [2:0] v3_1584201168_369;
   wire [2:0] v3_1584201168_370;
   wire [2:0] v3_1584201168_371;
   wire [2:0] v3_1584201168_372;
   wire [2:0] v3_1584201168_373;
   wire [2:0] v3_1584201168_374;
   wire [2:0] v3_1584201168_375;
   wire [2:0] v3_1584201168_376;
   wire [2:0] v3_1584201168_377;
   wire [2:0] v3_1584201168_378;
   wire v3_1584201168_379;
   wire [3:0] v3_1584201168_380;
   wire [3:0] v3_1584201168_381;
   wire [3:0] v3_1584201168_382;
   wire [3:0] v3_1584201168_383;
   wire [3:0] v3_1584201168_384;
   wire [3:0] v3_1584201168_385;
   wire [2:0] v3_1584201168_386;
   wire [2:0] v3_1584201168_387;
   wire [2:0] v3_1584201168_388;
   wire [2:0] v3_1584201168_389;
   wire [2:0] v3_1584201168_390;
   wire [2:0] v3_1584201168_391;
   wire [2:0] v3_1584201168_392;
   wire [2:0] v3_1584201168_393;
   wire [2:0] v3_1584201168_394;
   wire [2:0] v3_1584201168_395;
   wire [2:0] v3_1584201168_396;
   wire [2:0] v3_1584201168_397;
   wire [2:0] v3_1584201168_398;
   wire [2:0] v3_1584201168_399;
   wire [2:0] v3_1584201168_400;
   wire [2:0] v3_1584201168_401;
   wire [2:0] v3_1584201168_402;
   wire [2:0] v3_1584201168_403;
   wire [2:0] v3_1584201168_404;
   wire [2:0] v3_1584201168_405;
   wire [2:0] v3_1584201168_406;
   wire [2:0] v3_1584201168_407;
   wire [2:0] v3_1584201168_408;
   wire [2:0] v3_1584201168_409;
   wire [2:0] v3_1584201168_410;
   wire v3_1584201168_411;
   wire [3:0] v3_1584201168_412;
   wire [3:0] v3_1584201168_413;
   wire [3:0] v3_1584201168_414;
   wire [3:0] v3_1584201168_415;
   wire [3:0] v3_1584201168_416;
   wire [3:0] v3_1584201168_417;
   wire [2:0] v3_1584201168_418;
   wire [2:0] v3_1584201168_419;
   wire v3_1584201168_420;
   wire v3_1584201168_421;
   wire v3_1584201168_422;
   wire v3_1584201168_423;
   wire v3_1584201168_424;
   wire v3_1584201168_425;
   wire v3_1584201168_426;
   wire v3_1584201168_427;
   wire [7:0] v3_1584201168_428;
   wire [7:0] v3_1584201168_429;
   wire [7:0] v3_1584201168_430;
   wire [7:0] v3_1584201168_431;
   wire [7:0] v3_1584201168_432;
   wire [4:0] v3_1584201168_433;
   wire [7:0] v3_1584201168_434;
   wire [7:0] v3_1584201168_435;
   wire [7:0] v3_1584201168_436;
   wire [7:0] v3_1584201168_437;
   wire [7:0] v3_1584201168_438;
   wire [7:0] v3_1584201168_439;
   wire [7:0] v3_1584201168_440;
   wire [7:0] v3_1584201168_441;
   wire [7:0] v3_1584201168_442;
   wire [7:0] v3_1584201168_443;
   wire [7:0] v3_1584201168_444;
   wire [7:0] v3_1584201168_445;
   wire [7:0] v3_1584201168_446;
   wire [7:0] v3_1584201168_447;
   wire [7:0] v3_1584201168_448;
   wire [7:0] v3_1584201168_449;
   wire [7:0] v3_1584201168_450;
   wire v3_1584201168_451;

   // Output Net Declarations
   wire p;
   wire [2:0] coinOutNTD_50;
   wire [2:0] coinOutNTD_10;
   wire [2:0] coinOutNTD_5;
   wire [2:0] coinOutNTD_1;
   wire [1:0] itemTypeOut;
   wire [1:0] serviceTypeOut;

   // Combinational Assignments
   assign v3_1584201168_0 = 1'b0; 
   assign v3_1584201168_23 = v3_1584201168_62 ? v3_1584201168_61 : v3_1584201168_24;
   assign v3_1584201168_24 = v3_1584201168_25;
   assign v3_1584201168_25 = v3_1584201168_60 ? v3_1584201168_56 : v3_1584201168_26;
   assign v3_1584201168_26 = v3_1584201168_55 ? v3_1584201168_54 : v3_1584201168_27;
   assign v3_1584201168_27 = v3_1584201168_53 ? v3_1584201168_32 : v3_1584201168_28;
   assign v3_1584201168_28 = v3_1584201168_51 ? v3_1584201168_43 : v3_1584201168_29;
   assign v3_1584201168_29 = v3_1584201168_41 ? v3_1584201168_32 : v3_1584201168_30;
   assign v3_1584201168_30 = v3_1584201168_39 ? v3_1584201168_32 : v3_1584201168_31;
   assign v3_1584201168_31 = v3_1584201168_37 ? v3_1584201168_33 : v3_1584201168_32;
   assign v3_1584201168_32 = v3_1584201168_8;
   assign v3_1584201168_33 = v3_1584201168_36 ? v3_1584201168_34 : v3_1584201168_32;
   assign v3_1584201168_34 = v3_1584201168_35;
   assign v3_1584201168_35 = 3'b000; 
   assign v3_1584201168_36 = v3_1584201168_21 == v3_1584201168_35;
   assign v3_1584201168_37 = v3_1584201168_18 >= v3_1584201168_38;
   assign v3_1584201168_38 = 8'b00000001; 
   assign v3_1584201168_39 = v3_1584201168_17 == v3_1584201168_40;
   assign v3_1584201168_40 = 2'b10; 
   assign v3_1584201168_41 = v3_1584201168_17 == v3_1584201168_42;
   assign v3_1584201168_42 = 2'b01; 
   assign v3_1584201168_43 = v3_1584201168_49 ? v3_1584201168_44 : v3_1584201168_32;
   assign v3_1584201168_44 = v3_1584201168_48 ? v3_1584201168_32 : v3_1584201168_45;
   assign v3_1584201168_45 = v3_1584201168_47;
   assign v3_1584201168_46 = 3'b001; 
   assign v3_1584201168_47 = v3_1584201168_8 + v3_1584201168_46;
   assign v3_1584201168_48 = v3_1584201168_19 == v3_1584201168_35;
   assign v3_1584201168_49 = v3_1584201168_18 >= v3_1584201168_50;
   assign v3_1584201168_50 = 8'b00110010; 
   assign v3_1584201168_51 = v3_1584201168_17 == v3_1584201168_52;
   assign v3_1584201168_52 = 2'b00; 
   assign v3_1584201168_53 = ~v3_1584201168_16;
   assign v3_1584201168_54 = v3_1584201168_35;
   assign v3_1584201168_55 = v3_1584201168_13 == v3_1584201168_52;
   assign v3_1584201168_56 = v3_1584201168_58 ? v3_1584201168_57 : v3_1584201168_32;
   assign v3_1584201168_57 = v3_1584201168_35;
   assign v3_1584201168_58 = ~v3_1584201168_59;
   assign v3_1584201168_59 = itemTypeIn == v3_1584201168_52;
   assign v3_1584201168_60 = v3_1584201168_13 == v3_1584201168_42;
   assign v3_1584201168_61 = v3_1584201168_35;
   assign v3_1584201168_62 = ~reset;
   assign v3_1584201168_63 = 3'b000; 
   assign v3_1584201168_64 = v3_1584201168_62 ? v3_1584201168_86 : v3_1584201168_65;
   assign v3_1584201168_65 = v3_1584201168_66;
   assign v3_1584201168_66 = v3_1584201168_60 ? v3_1584201168_84 : v3_1584201168_67;
   assign v3_1584201168_67 = v3_1584201168_55 ? v3_1584201168_83 : v3_1584201168_68;
   assign v3_1584201168_68 = v3_1584201168_53 ? v3_1584201168_73 : v3_1584201168_69;
   assign v3_1584201168_69 = v3_1584201168_51 ? v3_1584201168_73 : v3_1584201168_70;
   assign v3_1584201168_70 = v3_1584201168_41 ? v3_1584201168_76 : v3_1584201168_71;
   assign v3_1584201168_71 = v3_1584201168_39 ? v3_1584201168_73 : v3_1584201168_72;
   assign v3_1584201168_72 = v3_1584201168_37 ? v3_1584201168_74 : v3_1584201168_73;
   assign v3_1584201168_73 = v3_1584201168_9;
   assign v3_1584201168_74 = v3_1584201168_36 ? v3_1584201168_75 : v3_1584201168_73;
   assign v3_1584201168_75 = v3_1584201168_35;
   assign v3_1584201168_76 = v3_1584201168_81 ? v3_1584201168_77 : v3_1584201168_73;
   assign v3_1584201168_77 = v3_1584201168_80 ? v3_1584201168_73 : v3_1584201168_78;
   assign v3_1584201168_78 = v3_1584201168_79;
   assign v3_1584201168_79 = v3_1584201168_9 + v3_1584201168_46;
   assign v3_1584201168_80 = v3_1584201168_20 == v3_1584201168_35;
   assign v3_1584201168_81 = v3_1584201168_18 >= v3_1584201168_82;
   assign v3_1584201168_82 = 8'b00001010; 
   assign v3_1584201168_83 = v3_1584201168_35;
   assign v3_1584201168_84 = v3_1584201168_58 ? v3_1584201168_85 : v3_1584201168_73;
   assign v3_1584201168_85 = v3_1584201168_35;
   assign v3_1584201168_86 = v3_1584201168_35;
   assign v3_1584201168_87 = 3'b000; 
   assign v3_1584201168_88 = v3_1584201168_62 ? v3_1584201168_110 : v3_1584201168_89;
   assign v3_1584201168_89 = v3_1584201168_90;
   assign v3_1584201168_90 = v3_1584201168_60 ? v3_1584201168_108 : v3_1584201168_91;
   assign v3_1584201168_91 = v3_1584201168_55 ? v3_1584201168_107 : v3_1584201168_92;
   assign v3_1584201168_92 = v3_1584201168_53 ? v3_1584201168_97 : v3_1584201168_93;
   assign v3_1584201168_93 = v3_1584201168_51 ? v3_1584201168_97 : v3_1584201168_94;
   assign v3_1584201168_94 = v3_1584201168_41 ? v3_1584201168_97 : v3_1584201168_95;
   assign v3_1584201168_95 = v3_1584201168_39 ? v3_1584201168_100 : v3_1584201168_96;
   assign v3_1584201168_96 = v3_1584201168_37 ? v3_1584201168_98 : v3_1584201168_97;
   assign v3_1584201168_97 = v3_1584201168_10;
   assign v3_1584201168_98 = v3_1584201168_36 ? v3_1584201168_99 : v3_1584201168_97;
   assign v3_1584201168_99 = v3_1584201168_35;
   assign v3_1584201168_100 = v3_1584201168_105 ? v3_1584201168_101 : v3_1584201168_97;
   assign v3_1584201168_101 = v3_1584201168_104 ? v3_1584201168_97 : v3_1584201168_102;
   assign v3_1584201168_102 = v3_1584201168_103;
   assign v3_1584201168_103 = v3_1584201168_10 + v3_1584201168_46;
   assign v3_1584201168_104 = v3_1584201168_22 == v3_1584201168_35;
   assign v3_1584201168_105 = v3_1584201168_18 >= v3_1584201168_106;
   assign v3_1584201168_106 = 8'b00000101; 
   assign v3_1584201168_107 = v3_1584201168_35;
   assign v3_1584201168_108 = v3_1584201168_58 ? v3_1584201168_109 : v3_1584201168_97;
   assign v3_1584201168_109 = v3_1584201168_35;
   assign v3_1584201168_110 = v3_1584201168_35;
   assign v3_1584201168_111 = 3'b000; 
   assign v3_1584201168_112 = v3_1584201168_62 ? v3_1584201168_129 : v3_1584201168_113;
   assign v3_1584201168_113 = v3_1584201168_114;
   assign v3_1584201168_114 = v3_1584201168_60 ? v3_1584201168_127 : v3_1584201168_115;
   assign v3_1584201168_115 = v3_1584201168_55 ? v3_1584201168_126 : v3_1584201168_116;
   assign v3_1584201168_116 = v3_1584201168_53 ? v3_1584201168_121 : v3_1584201168_117;
   assign v3_1584201168_117 = v3_1584201168_51 ? v3_1584201168_121 : v3_1584201168_118;
   assign v3_1584201168_118 = v3_1584201168_41 ? v3_1584201168_121 : v3_1584201168_119;
   assign v3_1584201168_119 = v3_1584201168_39 ? v3_1584201168_121 : v3_1584201168_120;
   assign v3_1584201168_120 = v3_1584201168_37 ? v3_1584201168_122 : v3_1584201168_121;
   assign v3_1584201168_121 = v3_1584201168_11;
   assign v3_1584201168_122 = v3_1584201168_36 ? v3_1584201168_125 : v3_1584201168_123;
   assign v3_1584201168_123 = v3_1584201168_124;
   assign v3_1584201168_124 = v3_1584201168_11 + v3_1584201168_46;
   assign v3_1584201168_125 = v3_1584201168_35;
   assign v3_1584201168_126 = v3_1584201168_35;
   assign v3_1584201168_127 = v3_1584201168_58 ? v3_1584201168_128 : v3_1584201168_121;
   assign v3_1584201168_128 = v3_1584201168_35;
   assign v3_1584201168_129 = v3_1584201168_35;
   assign v3_1584201168_130 = 3'b000; 
   assign v3_1584201168_131 = v3_1584201168_62 ? v3_1584201168_150 : v3_1584201168_132;
   assign v3_1584201168_132 = v3_1584201168_133;
   assign v3_1584201168_133 = v3_1584201168_60 ? v3_1584201168_148 : v3_1584201168_134;
   assign v3_1584201168_134 = v3_1584201168_55 ? v3_1584201168_147 : v3_1584201168_135;
   assign v3_1584201168_135 = v3_1584201168_53 ? v3_1584201168_143 : v3_1584201168_136;
   assign v3_1584201168_136 = v3_1584201168_51 ? v3_1584201168_140 : v3_1584201168_137;
   assign v3_1584201168_137 = v3_1584201168_41 ? v3_1584201168_140 : v3_1584201168_138;
   assign v3_1584201168_138 = v3_1584201168_39 ? v3_1584201168_140 : v3_1584201168_139;
   assign v3_1584201168_139 = v3_1584201168_37 ? v3_1584201168_141 : v3_1584201168_140;
   assign v3_1584201168_140 = v3_1584201168_12;
   assign v3_1584201168_141 = v3_1584201168_36 ? v3_1584201168_142 : v3_1584201168_140;
   assign v3_1584201168_142 = v3_1584201168_52;
   assign v3_1584201168_143 = v3_1584201168_145 ? v3_1584201168_144 : v3_1584201168_140;
   assign v3_1584201168_144 = v3_1584201168_52;
   assign v3_1584201168_145 = ~v3_1584201168_146;
   assign v3_1584201168_146 = v3_1584201168_15 >= v3_1584201168_18;
   assign v3_1584201168_147 = v3_1584201168_52;
   assign v3_1584201168_148 = v3_1584201168_58 ? v3_1584201168_149 : v3_1584201168_140;
   assign v3_1584201168_149 = itemTypeIn;
   assign v3_1584201168_150 = v3_1584201168_52;
   assign v3_1584201168_151 = 2'b00; 
   assign v3_1584201168_152 = v3_1584201168_62 ? v3_1584201168_168 : v3_1584201168_153;
   assign v3_1584201168_153 = v3_1584201168_154;
   assign v3_1584201168_154 = v3_1584201168_60 ? v3_1584201168_166 : v3_1584201168_155;
   assign v3_1584201168_155 = v3_1584201168_55 ? v3_1584201168_165 : v3_1584201168_156;
   assign v3_1584201168_156 = v3_1584201168_53 ? v3_1584201168_163 : v3_1584201168_157;
   assign v3_1584201168_157 = v3_1584201168_51 ? v3_1584201168_163 : v3_1584201168_158;
   assign v3_1584201168_158 = v3_1584201168_41 ? v3_1584201168_163 : v3_1584201168_159;
   assign v3_1584201168_159 = v3_1584201168_39 ? v3_1584201168_163 : v3_1584201168_160;
   assign v3_1584201168_160 = v3_1584201168_37 ? v3_1584201168_162 : v3_1584201168_161;
   assign v3_1584201168_161 = v3_1584201168_52;
   assign v3_1584201168_162 = v3_1584201168_36 ? v3_1584201168_164 : v3_1584201168_163;
   assign v3_1584201168_163 = v3_1584201168_13;
   assign v3_1584201168_164 = v3_1584201168_52;
   assign v3_1584201168_165 = v3_1584201168_42;
   assign v3_1584201168_166 = v3_1584201168_58 ? v3_1584201168_167 : v3_1584201168_163;
   assign v3_1584201168_167 = v3_1584201168_40;
   assign v3_1584201168_168 = v3_1584201168_42;
   assign v3_1584201168_169 = 2'b00; 
   assign v3_1584201168_170 = v3_1584201168_62 ? v3_1584201168_172 : v3_1584201168_171;
   assign v3_1584201168_171 = v3_1584201168_14;
   assign v3_1584201168_172 = v3_1584201168_173;
   assign v3_1584201168_173 = 1'b1; 
   assign v3_1584201168_174 = 1'b0; 
   assign v3_1584201168_175 = v3_1584201168_62 ? v3_1584201168_203 : v3_1584201168_176;
   assign v3_1584201168_176 = v3_1584201168_177;
   assign v3_1584201168_177 = v3_1584201168_60 ? v3_1584201168_179 : v3_1584201168_178;
   assign v3_1584201168_178 = v3_1584201168_15;
   assign v3_1584201168_179 = v3_1584201168_58 ? v3_1584201168_180 : v3_1584201168_178;
   assign v3_1584201168_180 = v3_1584201168_202;
   assign v3_1584201168_181 = v3_1584201168_197;
   assign v3_1584201168_182 = v3_1584201168_192;
   assign v3_1584201168_183 = v3_1584201168_187;
   assign v3_1584201168_184 = v3_1584201168_186;
   assign v3_1584201168_185 = 6'b000000; 
   assign v3_1584201168_186 = {v3_1584201168_185, coinInNTD_50};
   assign v3_1584201168_187 = v3_1584201168_50 * v3_1584201168_184;
   assign v3_1584201168_188 = v3_1584201168_191;
   assign v3_1584201168_189 = v3_1584201168_190;
   assign v3_1584201168_190 = {v3_1584201168_185, coinInNTD_10};
   assign v3_1584201168_191 = v3_1584201168_82 * v3_1584201168_189;
   assign v3_1584201168_192 = v3_1584201168_183 + v3_1584201168_188;
   assign v3_1584201168_193 = v3_1584201168_196;
   assign v3_1584201168_194 = v3_1584201168_195;
   assign v3_1584201168_195 = {v3_1584201168_185, coinInNTD_5};
   assign v3_1584201168_196 = v3_1584201168_106 * v3_1584201168_194;
   assign v3_1584201168_197 = v3_1584201168_182 + v3_1584201168_193;
   assign v3_1584201168_198 = v3_1584201168_201;
   assign v3_1584201168_199 = v3_1584201168_200;
   assign v3_1584201168_200 = {v3_1584201168_185, coinInNTD_1};
   assign v3_1584201168_201 = v3_1584201168_38 * v3_1584201168_199;
   assign v3_1584201168_202 = v3_1584201168_181 + v3_1584201168_198;
   assign v3_1584201168_203 = v3_1584201168_204;
   assign v3_1584201168_204 = 8'b00000000; 
   assign v3_1584201168_205 = 8'b00000000; 
   assign v3_1584201168_206 = v3_1584201168_62 ? v3_1584201168_218 : v3_1584201168_207;
   assign v3_1584201168_207 = v3_1584201168_208;
   assign v3_1584201168_208 = v3_1584201168_60 ? v3_1584201168_215 : v3_1584201168_209;
   assign v3_1584201168_209 = v3_1584201168_55 ? v3_1584201168_211 : v3_1584201168_210;
   assign v3_1584201168_210 = v3_1584201168_53 ? v3_1584201168_212 : v3_1584201168_211;
   assign v3_1584201168_211 = v3_1584201168_16;
   assign v3_1584201168_212 = v3_1584201168_145 ? v3_1584201168_214 : v3_1584201168_213;
   assign v3_1584201168_213 = v3_1584201168_173;
   assign v3_1584201168_214 = v3_1584201168_173;
   assign v3_1584201168_215 = v3_1584201168_58 ? v3_1584201168_216 : v3_1584201168_211;
   assign v3_1584201168_216 = v3_1584201168_217;
   assign v3_1584201168_217 = 1'b0; 
   assign v3_1584201168_218 = v3_1584201168_217;
   assign v3_1584201168_219 = 1'b0; 
   assign v3_1584201168_220 = v3_1584201168_62 ? v3_1584201168_247 : v3_1584201168_221;
   assign v3_1584201168_221 = v3_1584201168_222;
   assign v3_1584201168_222 = v3_1584201168_60 ? v3_1584201168_245 : v3_1584201168_223;
   assign v3_1584201168_223 = v3_1584201168_55 ? v3_1584201168_229 : v3_1584201168_224;
   assign v3_1584201168_224 = v3_1584201168_53 ? v3_1584201168_229 : v3_1584201168_225;
   assign v3_1584201168_225 = v3_1584201168_51 ? v3_1584201168_241 : v3_1584201168_226;
   assign v3_1584201168_226 = v3_1584201168_41 ? v3_1584201168_237 : v3_1584201168_227;
   assign v3_1584201168_227 = v3_1584201168_39 ? v3_1584201168_232 : v3_1584201168_228;
   assign v3_1584201168_228 = v3_1584201168_37 ? v3_1584201168_230 : v3_1584201168_229;
   assign v3_1584201168_229 = v3_1584201168_17;
   assign v3_1584201168_230 = v3_1584201168_36 ? v3_1584201168_231 : v3_1584201168_229;
   assign v3_1584201168_231 = v3_1584201168_52;
   assign v3_1584201168_232 = v3_1584201168_105 ? v3_1584201168_235 : v3_1584201168_233;
   assign v3_1584201168_233 = v3_1584201168_234;
   assign v3_1584201168_234 = 2'b11; 
   assign v3_1584201168_235 = v3_1584201168_104 ? v3_1584201168_236 : v3_1584201168_229;
   assign v3_1584201168_236 = v3_1584201168_234;
   assign v3_1584201168_237 = v3_1584201168_81 ? v3_1584201168_239 : v3_1584201168_238;
   assign v3_1584201168_238 = v3_1584201168_40;
   assign v3_1584201168_239 = v3_1584201168_80 ? v3_1584201168_240 : v3_1584201168_229;
   assign v3_1584201168_240 = v3_1584201168_40;
   assign v3_1584201168_241 = v3_1584201168_49 ? v3_1584201168_243 : v3_1584201168_242;
   assign v3_1584201168_242 = v3_1584201168_42;
   assign v3_1584201168_243 = v3_1584201168_48 ? v3_1584201168_244 : v3_1584201168_229;
   assign v3_1584201168_244 = v3_1584201168_42;
   assign v3_1584201168_245 = v3_1584201168_58 ? v3_1584201168_246 : v3_1584201168_229;
   assign v3_1584201168_246 = v3_1584201168_52;
   assign v3_1584201168_247 = v3_1584201168_52;
   assign v3_1584201168_248 = 2'b00; 
   assign v3_1584201168_249 = v3_1584201168_62 ? v3_1584201168_289 : v3_1584201168_250;
   assign v3_1584201168_250 = v3_1584201168_251;
   assign v3_1584201168_251 = v3_1584201168_60 ? v3_1584201168_279 : v3_1584201168_252;
   assign v3_1584201168_252 = v3_1584201168_55 ? v3_1584201168_258 : v3_1584201168_253;
   assign v3_1584201168_253 = v3_1584201168_53 ? v3_1584201168_275 : v3_1584201168_254;
   assign v3_1584201168_254 = v3_1584201168_51 ? v3_1584201168_271 : v3_1584201168_255;
   assign v3_1584201168_255 = v3_1584201168_41 ? v3_1584201168_267 : v3_1584201168_256;
   assign v3_1584201168_256 = v3_1584201168_39 ? v3_1584201168_263 : v3_1584201168_257;
   assign v3_1584201168_257 = v3_1584201168_37 ? v3_1584201168_259 : v3_1584201168_258;
   assign v3_1584201168_258 = v3_1584201168_18;
   assign v3_1584201168_259 = v3_1584201168_36 ? v3_1584201168_262 : v3_1584201168_260;
   assign v3_1584201168_260 = v3_1584201168_261;
   assign v3_1584201168_261 = v3_1584201168_18 - v3_1584201168_38;
   assign v3_1584201168_262 = v3_1584201168_15;
   assign v3_1584201168_263 = v3_1584201168_105 ? v3_1584201168_264 : v3_1584201168_258;
   assign v3_1584201168_264 = v3_1584201168_104 ? v3_1584201168_258 : v3_1584201168_265;
   assign v3_1584201168_265 = v3_1584201168_266;
   assign v3_1584201168_266 = v3_1584201168_18 - v3_1584201168_106;
   assign v3_1584201168_267 = v3_1584201168_81 ? v3_1584201168_268 : v3_1584201168_258;
   assign v3_1584201168_268 = v3_1584201168_80 ? v3_1584201168_258 : v3_1584201168_269;
   assign v3_1584201168_269 = v3_1584201168_270;
   assign v3_1584201168_270 = v3_1584201168_18 - v3_1584201168_82;
   assign v3_1584201168_271 = v3_1584201168_49 ? v3_1584201168_272 : v3_1584201168_258;
   assign v3_1584201168_272 = v3_1584201168_48 ? v3_1584201168_258 : v3_1584201168_273;
   assign v3_1584201168_273 = v3_1584201168_274;
   assign v3_1584201168_274 = v3_1584201168_18 - v3_1584201168_50;
   assign v3_1584201168_275 = v3_1584201168_145 ? v3_1584201168_278 : v3_1584201168_276;
   assign v3_1584201168_276 = v3_1584201168_277;
   assign v3_1584201168_277 = v3_1584201168_15 - v3_1584201168_18;
   assign v3_1584201168_278 = v3_1584201168_15;
   assign v3_1584201168_279 = v3_1584201168_58 ? v3_1584201168_280 : v3_1584201168_258;
   assign v3_1584201168_280 = v3_1584201168_288 ? v3_1584201168_287 : v3_1584201168_281;
   assign v3_1584201168_281 = v3_1584201168_286 ? v3_1584201168_285 : v3_1584201168_282;
   assign v3_1584201168_282 = v3_1584201168_284 ? v3_1584201168_283 : v3_1584201168_204;
   assign v3_1584201168_283 = 8'b00010110; 
   assign v3_1584201168_284 = itemTypeIn == v3_1584201168_234;
   assign v3_1584201168_285 = 8'b00001111; 
   assign v3_1584201168_286 = itemTypeIn == v3_1584201168_40;
   assign v3_1584201168_287 = 8'b00001000; 
   assign v3_1584201168_288 = itemTypeIn == v3_1584201168_42;
   assign v3_1584201168_289 = v3_1584201168_204;
   assign v3_1584201168_290 = 8'b00000000; 
   assign v3_1584201168_291 = v3_1584201168_62 ? v3_1584201168_323 : v3_1584201168_292;
   assign v3_1584201168_292 = v3_1584201168_293;
   assign v3_1584201168_293 = v3_1584201168_60 ? v3_1584201168_308 : v3_1584201168_294;
   assign v3_1584201168_294 = v3_1584201168_55 ? v3_1584201168_300 : v3_1584201168_295;
   assign v3_1584201168_295 = v3_1584201168_53 ? v3_1584201168_300 : v3_1584201168_296;
   assign v3_1584201168_296 = v3_1584201168_51 ? v3_1584201168_304 : v3_1584201168_297;
   assign v3_1584201168_297 = v3_1584201168_41 ? v3_1584201168_300 : v3_1584201168_298;
   assign v3_1584201168_298 = v3_1584201168_39 ? v3_1584201168_300 : v3_1584201168_299;
   assign v3_1584201168_299 = v3_1584201168_37 ? v3_1584201168_301 : v3_1584201168_300;
   assign v3_1584201168_300 = v3_1584201168_19;
   assign v3_1584201168_301 = v3_1584201168_36 ? v3_1584201168_302 : v3_1584201168_300;
   assign v3_1584201168_302 = v3_1584201168_303;
   assign v3_1584201168_303 = v3_1584201168_19 + v3_1584201168_8;
   assign v3_1584201168_304 = v3_1584201168_49 ? v3_1584201168_305 : v3_1584201168_300;
   assign v3_1584201168_305 = v3_1584201168_48 ? v3_1584201168_300 : v3_1584201168_306;
   assign v3_1584201168_306 = v3_1584201168_307;
   assign v3_1584201168_307 = v3_1584201168_19 - v3_1584201168_46;
   assign v3_1584201168_308 = v3_1584201168_58 ? v3_1584201168_309 : v3_1584201168_300;
   assign v3_1584201168_309 = v3_1584201168_315 ? v3_1584201168_314 : v3_1584201168_310;
   assign v3_1584201168_310 = v3_1584201168_313;
   assign v3_1584201168_311 = v3_1584201168_312;
   assign v3_1584201168_312 = {v3_1584201168_217, coinInNTD_50};
   assign v3_1584201168_313 = v3_1584201168_19 + v3_1584201168_311;
   assign v3_1584201168_314 = 3'b111; 
   assign v3_1584201168_315 = v3_1584201168_316 >= v3_1584201168_322;
   assign v3_1584201168_316 = v3_1584201168_321;
   assign v3_1584201168_317 = v3_1584201168_318;
   assign v3_1584201168_318 = {v3_1584201168_217, v3_1584201168_19};
   assign v3_1584201168_319 = v3_1584201168_320;
   assign v3_1584201168_320 = {v3_1584201168_52, coinInNTD_50};
   assign v3_1584201168_321 = v3_1584201168_317 + v3_1584201168_319;
   assign v3_1584201168_322 = 4'b0111; 
   assign v3_1584201168_323 = v3_1584201168_324;
   assign v3_1584201168_324 = 3'b010; 
   assign v3_1584201168_325 = 3'b000; 
   assign v3_1584201168_326 = v3_1584201168_62 ? v3_1584201168_356 : v3_1584201168_327;
   assign v3_1584201168_327 = v3_1584201168_328;
   assign v3_1584201168_328 = v3_1584201168_60 ? v3_1584201168_343 : v3_1584201168_329;
   assign v3_1584201168_329 = v3_1584201168_55 ? v3_1584201168_335 : v3_1584201168_330;
   assign v3_1584201168_330 = v3_1584201168_53 ? v3_1584201168_335 : v3_1584201168_331;
   assign v3_1584201168_331 = v3_1584201168_51 ? v3_1584201168_335 : v3_1584201168_332;
   assign v3_1584201168_332 = v3_1584201168_41 ? v3_1584201168_339 : v3_1584201168_333;
   assign v3_1584201168_333 = v3_1584201168_39 ? v3_1584201168_335 : v3_1584201168_334;
   assign v3_1584201168_334 = v3_1584201168_37 ? v3_1584201168_336 : v3_1584201168_335;
   assign v3_1584201168_335 = v3_1584201168_20;
   assign v3_1584201168_336 = v3_1584201168_36 ? v3_1584201168_337 : v3_1584201168_335;
   assign v3_1584201168_337 = v3_1584201168_338;
   assign v3_1584201168_338 = v3_1584201168_20 + v3_1584201168_9;
   assign v3_1584201168_339 = v3_1584201168_81 ? v3_1584201168_340 : v3_1584201168_335;
   assign v3_1584201168_340 = v3_1584201168_80 ? v3_1584201168_335 : v3_1584201168_341;
   assign v3_1584201168_341 = v3_1584201168_342;
   assign v3_1584201168_342 = v3_1584201168_20 - v3_1584201168_46;
   assign v3_1584201168_343 = v3_1584201168_58 ? v3_1584201168_344 : v3_1584201168_335;
   assign v3_1584201168_344 = v3_1584201168_349 ? v3_1584201168_314 : v3_1584201168_345;
   assign v3_1584201168_345 = v3_1584201168_348;
   assign v3_1584201168_346 = v3_1584201168_347;
   assign v3_1584201168_347 = {v3_1584201168_217, coinInNTD_10};
   assign v3_1584201168_348 = v3_1584201168_20 + v3_1584201168_346;
   assign v3_1584201168_349 = v3_1584201168_350 >= v3_1584201168_322;
   assign v3_1584201168_350 = v3_1584201168_355;
   assign v3_1584201168_351 = v3_1584201168_352;
   assign v3_1584201168_352 = {v3_1584201168_217, v3_1584201168_20};
   assign v3_1584201168_353 = v3_1584201168_354;
   assign v3_1584201168_354 = {v3_1584201168_52, coinInNTD_10};
   assign v3_1584201168_355 = v3_1584201168_351 + v3_1584201168_353;
   assign v3_1584201168_356 = v3_1584201168_324;
   assign v3_1584201168_357 = 3'b000; 
   assign v3_1584201168_358 = v3_1584201168_62 ? v3_1584201168_386 : v3_1584201168_359;
   assign v3_1584201168_359 = v3_1584201168_360;
   assign v3_1584201168_360 = v3_1584201168_60 ? v3_1584201168_373 : v3_1584201168_361;
   assign v3_1584201168_361 = v3_1584201168_55 ? v3_1584201168_367 : v3_1584201168_362;
   assign v3_1584201168_362 = v3_1584201168_53 ? v3_1584201168_367 : v3_1584201168_363;
   assign v3_1584201168_363 = v3_1584201168_51 ? v3_1584201168_367 : v3_1584201168_364;
   assign v3_1584201168_364 = v3_1584201168_41 ? v3_1584201168_367 : v3_1584201168_365;
   assign v3_1584201168_365 = v3_1584201168_39 ? v3_1584201168_367 : v3_1584201168_366;
   assign v3_1584201168_366 = v3_1584201168_37 ? v3_1584201168_368 : v3_1584201168_367;
   assign v3_1584201168_367 = v3_1584201168_21;
   assign v3_1584201168_368 = v3_1584201168_36 ? v3_1584201168_371 : v3_1584201168_369;
   assign v3_1584201168_369 = v3_1584201168_370;
   assign v3_1584201168_370 = v3_1584201168_21 - v3_1584201168_46;
   assign v3_1584201168_371 = v3_1584201168_372;
   assign v3_1584201168_372 = v3_1584201168_21 + v3_1584201168_11;
   assign v3_1584201168_373 = v3_1584201168_58 ? v3_1584201168_374 : v3_1584201168_367;
   assign v3_1584201168_374 = v3_1584201168_379 ? v3_1584201168_314 : v3_1584201168_375;
   assign v3_1584201168_375 = v3_1584201168_378;
   assign v3_1584201168_376 = v3_1584201168_377;
   assign v3_1584201168_377 = {v3_1584201168_217, coinInNTD_1};
   assign v3_1584201168_378 = v3_1584201168_21 + v3_1584201168_376;
   assign v3_1584201168_379 = v3_1584201168_380 >= v3_1584201168_322;
   assign v3_1584201168_380 = v3_1584201168_385;
   assign v3_1584201168_381 = v3_1584201168_382;
   assign v3_1584201168_382 = {v3_1584201168_217, v3_1584201168_21};
   assign v3_1584201168_383 = v3_1584201168_384;
   assign v3_1584201168_384 = {v3_1584201168_52, coinInNTD_1};
   assign v3_1584201168_385 = v3_1584201168_381 + v3_1584201168_383;
   assign v3_1584201168_386 = v3_1584201168_324;
   assign v3_1584201168_387 = 3'b000; 
   assign v3_1584201168_388 = v3_1584201168_62 ? v3_1584201168_418 : v3_1584201168_389;
   assign v3_1584201168_389 = v3_1584201168_390;
   assign v3_1584201168_390 = v3_1584201168_60 ? v3_1584201168_405 : v3_1584201168_391;
   assign v3_1584201168_391 = v3_1584201168_55 ? v3_1584201168_397 : v3_1584201168_392;
   assign v3_1584201168_392 = v3_1584201168_53 ? v3_1584201168_397 : v3_1584201168_393;
   assign v3_1584201168_393 = v3_1584201168_51 ? v3_1584201168_397 : v3_1584201168_394;
   assign v3_1584201168_394 = v3_1584201168_41 ? v3_1584201168_397 : v3_1584201168_395;
   assign v3_1584201168_395 = v3_1584201168_39 ? v3_1584201168_401 : v3_1584201168_396;
   assign v3_1584201168_396 = v3_1584201168_37 ? v3_1584201168_398 : v3_1584201168_397;
   assign v3_1584201168_397 = v3_1584201168_22;
   assign v3_1584201168_398 = v3_1584201168_36 ? v3_1584201168_399 : v3_1584201168_397;
   assign v3_1584201168_399 = v3_1584201168_400;
   assign v3_1584201168_400 = v3_1584201168_22 + v3_1584201168_10;
   assign v3_1584201168_401 = v3_1584201168_105 ? v3_1584201168_402 : v3_1584201168_397;
   assign v3_1584201168_402 = v3_1584201168_104 ? v3_1584201168_397 : v3_1584201168_403;
   assign v3_1584201168_403 = v3_1584201168_404;
   assign v3_1584201168_404 = v3_1584201168_22 - v3_1584201168_46;
   assign v3_1584201168_405 = v3_1584201168_58 ? v3_1584201168_406 : v3_1584201168_397;
   assign v3_1584201168_406 = v3_1584201168_411 ? v3_1584201168_314 : v3_1584201168_407;
   assign v3_1584201168_407 = v3_1584201168_410;
   assign v3_1584201168_408 = v3_1584201168_409;
   assign v3_1584201168_409 = {v3_1584201168_217, coinInNTD_5};
   assign v3_1584201168_410 = v3_1584201168_22 + v3_1584201168_408;
   assign v3_1584201168_411 = v3_1584201168_412 >= v3_1584201168_322;
   assign v3_1584201168_412 = v3_1584201168_417;
   assign v3_1584201168_413 = v3_1584201168_414;
   assign v3_1584201168_414 = {v3_1584201168_217, v3_1584201168_22};
   assign v3_1584201168_415 = v3_1584201168_416;
   assign v3_1584201168_416 = {v3_1584201168_52, coinInNTD_5};
   assign v3_1584201168_417 = v3_1584201168_413 + v3_1584201168_415;
   assign v3_1584201168_418 = v3_1584201168_324;
   assign v3_1584201168_419 = 3'b000; 
   assign v3_1584201168_420 = v3_1584201168_451;
   assign v3_1584201168_421 = v3_1584201168_425;
   assign v3_1584201168_422 = v3_1584201168_423;
   assign v3_1584201168_423 = v3_1584201168_14 & v3_1584201168_55;
   assign v3_1584201168_424 = v3_1584201168_12 == v3_1584201168_52;
   assign v3_1584201168_425 = v3_1584201168_422 & v3_1584201168_424;
   assign v3_1584201168_426 = ~v3_1584201168_427;
   assign v3_1584201168_427 = v3_1584201168_428 == v3_1584201168_15;
   assign v3_1584201168_428 = v3_1584201168_450;
   assign v3_1584201168_429 = v3_1584201168_445;
   assign v3_1584201168_430 = v3_1584201168_440;
   assign v3_1584201168_431 = v3_1584201168_435;
   assign v3_1584201168_432 = v3_1584201168_434;
   assign v3_1584201168_433 = 5'b00000; 
   assign v3_1584201168_434 = {v3_1584201168_433, v3_1584201168_8};
   assign v3_1584201168_435 = v3_1584201168_50 * v3_1584201168_432;
   assign v3_1584201168_436 = v3_1584201168_439;
   assign v3_1584201168_437 = v3_1584201168_438;
   assign v3_1584201168_438 = {v3_1584201168_433, v3_1584201168_9};
   assign v3_1584201168_439 = v3_1584201168_82 * v3_1584201168_437;
   assign v3_1584201168_440 = v3_1584201168_431 + v3_1584201168_436;
   assign v3_1584201168_441 = v3_1584201168_444;
   assign v3_1584201168_442 = v3_1584201168_443;
   assign v3_1584201168_443 = {v3_1584201168_433, v3_1584201168_10};
   assign v3_1584201168_444 = v3_1584201168_106 * v3_1584201168_442;
   assign v3_1584201168_445 = v3_1584201168_430 + v3_1584201168_441;
   assign v3_1584201168_446 = v3_1584201168_449;
   assign v3_1584201168_447 = v3_1584201168_448;
   assign v3_1584201168_448 = {v3_1584201168_433, v3_1584201168_11};
   assign v3_1584201168_449 = v3_1584201168_38 * v3_1584201168_447;
   assign v3_1584201168_450 = v3_1584201168_429 + v3_1584201168_446;
   assign v3_1584201168_451 = v3_1584201168_421 & v3_1584201168_426;

   // Output Net Assignments
   assign p = v3_1584201168_420;
   assign coinOutNTD_50 = v3_1584201168_8;
   assign coinOutNTD_10 = v3_1584201168_9;
   assign coinOutNTD_5 = v3_1584201168_10;
   assign coinOutNTD_1 = v3_1584201168_11;
   assign itemTypeOut = v3_1584201168_12;
   assign serviceTypeOut = v3_1584201168_13;

   // Non-blocking Assignments
   always @ (posedge clk) begin
      v3_1584201168_8 <= v3_1584201168_23;
      v3_1584201168_9 <= v3_1584201168_64;
      v3_1584201168_10 <= v3_1584201168_88;
      v3_1584201168_11 <= v3_1584201168_112;
      v3_1584201168_12 <= v3_1584201168_131;
      v3_1584201168_13 <= v3_1584201168_152;
      v3_1584201168_14 <= v3_1584201168_170;
      v3_1584201168_15 <= v3_1584201168_175;
      v3_1584201168_16 <= v3_1584201168_206;
      v3_1584201168_17 <= v3_1584201168_220;
      v3_1584201168_18 <= v3_1584201168_249;
      v3_1584201168_19 <= v3_1584201168_291;
      v3_1584201168_20 <= v3_1584201168_326;
      v3_1584201168_21 <= v3_1584201168_358;
      v3_1584201168_22 <= v3_1584201168_388;
   end
endmodule
